//Author: Kai Hughes | 2026 
//SHA-256 Core Testbench for DUT
//Tests with NIST vectors and the Bitcoin genesis block

`timescale 1ns/1ps

module sha256_core_tb;

    logic clk;
    logic rst_n;
    
    logic start;
    logic [511:0] block_in;
    logic [255:0] hash_in;
    logic init_hash;
    logic busy;
    logic done;
    logic [255:0] hash_out;
    
    sha256_core dut (.*);
    
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end
    
    int test_num;
    int errors;
    logic [255:0] expected_hash;
    
    task reset_system();
        rst_n = 0;
        start = 0;
        block_in = '0;
        hash_in = '0;
        init_hash = 1;
        
        repeat(5) @(posedge clk);
        rst_n = 1;
        repeat(2) @(posedge clk);
        
        $display("[%0t] Reset complete", $time);
    endtask
    
    task sha256_hash(input logic [511:0] block, 
                     input logic [255:0] prev_hash,
                     input logic init);
        @(posedge clk);
        block_in = block;
        hash_in = prev_hash;
        init_hash = init;
        start = 1;
        
        @(posedge clk);
        start = 0;
        
        wait(done == 1);
        @(posedge clk);
        
        $display("[%0t] Hash complete", $time);
    endtask
    
    task check_result(input logic [255:0] expected, input string test_name);
        if (hash_out === expected) begin
            $display(" PASS: %s", test_name);
            $display("   Result: %064x", hash_out);
        end else begin
            $display(" FAIL: %s", test_name);
            $display("   Expected: %064x", expected);
            $display("   Got:      %064x", hash_out);
            errors++;
        end
        $display("");
    endtask
    
    initial begin
        $display("             ");
        $display("SHA-256 Core Test");
        $display("             \n");
        
        errors = 0;
        test_num = 0;
        
        reset_system();
        
        //test case 1
        test_num++;
        $display("Test %0d: Empty string", test_num);
        
        block_in = {8'h80, 504'h0};  // 0x80 followed by zeros
        block_in[63:0] = 64'h0;      // length field = 0
        
        expected_hash = 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855;
        
        sha256_hash(block_in, '0, 1'b1);
        check_result(expected_hash, "Empty string");
        
        // test case 2 
        test_num++;
        $display("Test %0d: Message 'abc'", test_num);
        
        // "abc" = 0x616263
        block_in = {24'h616263, 8'h80, 416'h0, 64'h0000000000000018};
        
        expected_hash = 256'hba7816bf8f01cfea414140de5dae2223b00361a396177a9cb410ff61f20015ad;
        
        sha256_hash(block_in, '0, 1'b1);
        check_result(expected_hash, "Message 'abc'");
        
        //test case 3 
        test_num++;
        $display("Test %0d: Double SHA-256 of 'hello'", test_num);
        
        //initial hash
        block_in = {40'h68656c6c6f, 8'h80, 400'h0, 64'h0000000000000028};
        
        sha256_hash(block_in, '0, 1'b1);
        $display("   First hash: %064x", hash_out);
        
        logic [255:0] temp;
        temp = hash_out;
        
        // hash 2 
        block_in = {temp, 8'h80, 184'h0, 64'h0000000000000100};
        
        sha256_hash(block_in, '0, 1'b1);
        $display("   Final hash: %064x", hash_out);
        
        expected_hash = 256'h9595c9df90075148eb06860365df33584b75bff782a510c6cd4883a419833d50;
        check_result(expected_hash, "Double SHA-256 of 'hello'");
        
        test_num++;
        $display("Test %0d: Bitcoin Genesis Block (Part 1)", test_num);
        
        logic [639:0] genesis_header;
        genesis_header = 640'h0100000000000000000000000000000000000000000000000000000000000000000000003ba3edfd7a7b12b27ac72c3e76768f617fc81bc3888a51323a9fb8aa4b1e5e4a29ab5f49ffff001d1dac2b7c;
        
        block_in = genesis_header[639:128];
        
        sha256_hash(block_in, '0, 1'b1);
        temp = hash_out;
        $display("   Block 0 done: %064x", hash_out);
        
        test_num++;
        $display("Test %0d: Bitcoin Genesis Block (Part 2)", test_num);
        
        //Last 16 bytes + padding
        block_in = {genesis_header[127:0], 8'h80, 312'h0, 64'h0000000000000280};
        
        sha256_hash(block_in, temp, 1'b0);
        temp = hash_out;
        $display("   Block 1 done (first SHA-256 complete): %064x", hash_out);
        
        test_num++;
        $display("Test %0d: Bitcoin Genesis Block (Second SHA-256)", test_num);
        
        //has the hash
        block_in = {temp, 8'h80, 184'h0, 64'h0000000000000100};
        
        sha256_hash(block_in, '0, 1'b1);
        
        // genesis block hash (big-endian)
        expected_hash = 256'h6fe28c0ab6f1b372c1a6a246ae63f74f931e8365e15a089c68d6190000000000;
        
        $display("   Final double SHA-256: %064x", hash_out);
        check_result(expected_hash, "Bitcoin Genesis Block");
        
        $display("   Bitcoin displays this in reverse byte order:");
        $display("   000000000019d6689c085ae165831e934ff763ae46a2a6c172b3f1b60a8ce26f");
        $display("");
        
        $display("             ");
        $display("Test Summary");
        $display("Total tests: %0d", test_num);
        $display("Errors: %0d", errors);
        
        if (errors == 0) begin
            $display("\nALL TESTS PASSED\n");
        end else begin
            $display("\n%0d TESTS FAILED\n", errors);
        end
        
        $display("             \n");
        
        #100;
        $finish;
    end
    
    // Dump waveforms
    initial begin
        $dumpfile("sha256_core_tb.vcd");
        $dumpvars(0, sha256_core_tb);
    end
    
    initial begin
        #1000000;
        $display("ERROR: Simulation timeout");
        $finish;
    end

endmodule